/users/student/mr111/hccheng22/private/pda/HW1/NangateOpenCellLibrary.lef